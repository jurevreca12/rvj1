// TBA..
