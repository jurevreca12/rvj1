// TBA¸
